module test(
	input key,
	output led
);

assign led = key;

endmodule
